library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDi : std_logic_vector(3 downto 0) := "1011";
  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin


  tmp(0) := "000" & x"4" & '0' & x"00";  --  LDI $0
  tmp(1) := "000" & x"5" & '0' & x"00";  --  STA $ZERO
  tmp(2) := "000" & x"0" & '0' & x"00";  --  
  tmp(3) := "000" & x"4" & '1' & x"FF";  --  LDI $511
  tmp(4) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
  tmp(5) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
  tmp(6) := "000" & x"0" & '0' & x"00";  --  
  tmp(7) := "000" & x"4" & '0' & x"00";  --  LDI $0
  tmp(8) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
  tmp(9) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
 tmp(10) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
 tmp(11) := "000" & x"5" & '1' & x"23";  --  STA $HEX3
 tmp(12) := "000" & x"5" & '1' & x"24";  --  STA $HEX4
 tmp(13) := "000" & x"5" & '1' & x"25";  --  STA $HEX5
 tmp(14) := "000" & x"0" & '0' & x"00";  --  
 tmp(15) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
 tmp(16) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
 tmp(17) := "000" & x"5" & '1' & x"01";  --  STA $LEDR8
 tmp(18) := "000" & x"0" & '0' & x"00";  --  
 tmp(19) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
 tmp(20) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
 tmp(21) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
 tmp(22) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
 tmp(23) := "000" & x"5" & '0' & x"06";  --  STA $DEZENA_MILHAR
 tmp(24) := "000" & x"5" & '0' & x"07";  --  STA $CENTENA_MILHAR
 tmp(25) := "000" & x"0" & '0' & x"00";  --  
 tmp(26) := "000" & x"4" & '0' & x"09";  --  LDI $9
 tmp(27) := "000" & x"5" & '0' & x"08";  --  STA $LIM_UNIDADE
 tmp(28) := "000" & x"5" & '0' & x"09";  --  STA $LIM_DEZENA
 tmp(29) := "000" & x"5" & '0' & x"0A";  --  STA $LIM_CENTENA
 tmp(30) := "000" & x"5" & '0' & x"0B";  --  STA $LIM_MILHAR
 tmp(31) := "000" & x"5" & '0' & x"0C";  --  STA $LIM_DEZENA_MILHAR
 tmp(32) := "000" & x"5" & '0' & x"0D";  --  STA $LIM_CENTENA_MILHAR
 tmp(33) := "000" & x"5" & '0' & x"0E";  --  STA $NOVE
 tmp(34) := "000" & x"0" & '0' & x"00";  --  
 tmp(35) := "000" & x"4" & '0' & x"01";  --  LDI $1
 tmp(36) := "000" & x"5" & '0' & x"0F";  --  STA $UM
 tmp(37) := "000" & x"0" & '0' & x"00";  --  
 tmp(38) := "000" & x"4" & '0' & x"02";  --  LDI $2
 tmp(39) := "000" & x"5" & '0' & x"10";  --  STA $DOIS
 tmp(40) := "000" & x"0" & '0' & x"00";  --  
 tmp(41) := "000" & x"4" & '0' & x"05";  --  LDI $5
 tmp(42) := "000" & x"5" & '0' & x"11";  --  STA $CINCO
 tmp(43) := "000" & x"0" & '0' & x"00";  --  
 tmp(44) := "000" & x"4" & '0' & x"03";  --  LDI $3
 tmp(45) := "000" & x"5" & '0' & x"12";  --  STA $TRES
 tmp(46) := "000" & x"0" & '0' & x"00";  --  
 tmp(47) := "000" & x"0" & '0' & x"00";  --  main_loop:
 tmp(48) := "000" & x"0" & '0' & x"00";  --  
 tmp(49) := "000" & x"1" & '1' & x"60";  --  LDA $KEY0
 tmp(50) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(51) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(52) := "000" & x"7" & '0' & x"36";  --  JEQ .nao_leu_key0
 tmp(53) := "000" & x"9" & '0' & x"A6";  --  JSR .incrementa
 tmp(54) := "000" & x"0" & '0' & x"00";  --  nao_leu_key0:
 tmp(55) := "000" & x"0" & '0' & x"00";  --  
 tmp(56) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
 tmp(57) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(58) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(59) := "000" & x"7" & '0' & x"3D";  --  JEQ .nao_leu_key1
 tmp(60) := "000" & x"9" & '0' & x"FD";  --  JSR .limite
 tmp(61) := "000" & x"0" & '0' & x"00";  --  nao_leu_key1:
 tmp(62) := "000" & x"0" & '0' & x"00";  --  
 tmp(63) := "000" & x"1" & '1' & x"64";  --  LDA $FPGA_RESET
 tmp(64) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(65) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(66) := "000" & x"7" & '0' & x"44";  --  JEQ .nao_reset
 tmp(67) := "000" & x"9" & '0' & x"99";  --  JSR .reset
 tmp(68) := "000" & x"0" & '0' & x"00";  --  nao_reset:
 tmp(69) := "000" & x"0" & '0' & x"00";  --  
 tmp(70) := "000" & x"9" & '0' & x"5C";  --  JSR .verifica_limite
 tmp(71) := "000" & x"0" & '0' & x"00";  --  
 tmp(72) := "000" & x"1" & '0' & x"02";  --  LDA $UNIDADE
 tmp(73) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
 tmp(74) := "000" & x"0" & '0' & x"00";  --  
 tmp(75) := "000" & x"1" & '0' & x"03";  --  LDA $DEZENA
 tmp(76) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
 tmp(77) := "000" & x"0" & '0' & x"00";  --  
 tmp(78) := "000" & x"1" & '0' & x"04";  --  LDA $CENTENA
 tmp(79) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
 tmp(80) := "000" & x"0" & '0' & x"00";  --  
 tmp(81) := "000" & x"1" & '0' & x"05";  --  LDA $MILHAR
 tmp(82) := "000" & x"5" & '1' & x"23";  --  STA $HEX3
 tmp(83) := "000" & x"0" & '0' & x"00";  --  
 tmp(84) := "000" & x"1" & '0' & x"06";  --  LDA $DEZENA_MILHAR
 tmp(85) := "000" & x"5" & '1' & x"24";  --  STA $HEX4
 tmp(86) := "000" & x"0" & '0' & x"00";  --  
 tmp(87) := "000" & x"1" & '0' & x"07";  --  LDA $CENTENA_MILHAR
 tmp(88) := "000" & x"5" & '1' & x"25";  --  STA $HEX5
 tmp(89) := "000" & x"0" & '0' & x"00";  --  
 tmp(90) := "000" & x"6" & '0' & x"2F";  --  JMP .main_loop
 tmp(91) := "000" & x"0" & '0' & x"00";  --  
 tmp(92) := "000" & x"0" & '0' & x"00";  --  verifica_limite:
 tmp(93) := "000" & x"0" & '0' & x"00";  --  verifica_unidade:
 tmp(94) := "000" & x"1" & '0' & x"02";  --  LDA $UNIDADE
 tmp(95) := "000" & x"8" & '0' & x"08";  --  CEQ $LIM_UNIDADE
 tmp(96) := "000" & x"7" & '0' & x"66";  --  JEQ .verifica_dezena
 tmp(97) := "000" & x"4" & '0' & x"00";  --  LDI $0
 tmp(98) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
 tmp(99) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(100) := "000" & x"A" & '0' & x"00";  --  RET
tmp(101) := "000" & x"0" & '0' & x"00";  --  
tmp(102) := "000" & x"0" & '0' & x"00";  --  verifica_dezena:
tmp(103) := "000" & x"1" & '0' & x"03";  --  LDA $DEZENA
tmp(104) := "000" & x"8" & '0' & x"09";  --  CEQ $LIM_DEZENA
tmp(105) := "000" & x"7" & '0' & x"6F";  --  JEQ .verifica_centena
tmp(106) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(107) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(108) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(109) := "000" & x"A" & '0' & x"00";  --  RET
tmp(110) := "000" & x"0" & '0' & x"00";  --  
tmp(111) := "000" & x"0" & '0' & x"00";  --  verifica_centena:
tmp(112) := "000" & x"1" & '0' & x"04";  --  LDA $CENTENA
tmp(113) := "000" & x"8" & '0' & x"0A";  --  CEQ $LIM_CENTENA
tmp(114) := "000" & x"7" & '0' & x"78";  --  JEQ .verifica_milhar
tmp(115) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(116) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(117) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(118) := "000" & x"A" & '0' & x"00";  --  RET
tmp(119) := "000" & x"0" & '0' & x"00";  --  
tmp(120) := "000" & x"0" & '0' & x"00";  --  verifica_milhar:
tmp(121) := "000" & x"1" & '0' & x"05";  --  LDA $MILHAR
tmp(122) := "000" & x"8" & '0' & x"0B";  --  CEQ $LIM_MILHAR
tmp(123) := "000" & x"7" & '0' & x"81";  --  JEQ .verifica_dezena_milhar
tmp(124) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(125) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(126) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(127) := "000" & x"A" & '0' & x"00";  --  RET
tmp(128) := "000" & x"0" & '0' & x"00";  --  
tmp(129) := "000" & x"0" & '0' & x"00";  --  verifica_dezena_milhar:
tmp(130) := "000" & x"1" & '0' & x"06";  --  LDA $DEZENA_MILHAR
tmp(131) := "000" & x"8" & '0' & x"0C";  --  CEQ $LIM_DEZENA_MILHAR
tmp(132) := "000" & x"7" & '0' & x"8A";  --  JEQ .verifica_centena_milhar
tmp(133) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(134) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(135) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(136) := "000" & x"A" & '0' & x"00";  --  RET
tmp(137) := "000" & x"0" & '0' & x"00";  --  
tmp(138) := "000" & x"0" & '0' & x"00";  --  verifica_centena_milhar:
tmp(139) := "000" & x"1" & '0' & x"07";  --  LDA $CENTENA_MILHAR
tmp(140) := "000" & x"8" & '0' & x"0D";  --  CEQ $LIM_CENTENA_MILHAR
tmp(141) := "000" & x"7" & '0' & x"93";  --  JEQ .habilita_flag
tmp(142) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(143) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(144) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(145) := "000" & x"A" & '0' & x"00";  --  RET
tmp(146) := "000" & x"0" & '0' & x"00";  --  
tmp(147) := "000" & x"0" & '0' & x"00";  --  habilita_flag:
tmp(148) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(149) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(150) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(151) := "000" & x"A" & '0' & x"00";  --  RET
tmp(152) := "000" & x"0" & '0' & x"00";  --  
tmp(153) := "000" & x"0" & '0' & x"00";  --  reset:
tmp(154) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(155) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(156) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(157) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(158) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
tmp(159) := "000" & x"5" & '0' & x"06";  --  STA $DEZENA_MILHAR
tmp(160) := "000" & x"5" & '0' & x"07";  --  STA $CENTENA_MILHAR
tmp(161) := "000" & x"5" & '0' & x"01";  --  STA $FLAG_INIBE_CONT
tmp(162) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
tmp(163) := "000" & x"5" & '1' & x"01";  --  STA $LEDR8
tmp(164) := "000" & x"A" & '0' & x"00";  --  RET
tmp(165) := "000" & x"0" & '0' & x"00";  --  
tmp(166) := "000" & x"0" & '0' & x"00";  --  incrementa:
tmp(167) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(168) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
tmp(169) := "000" & x"0" & '0' & x"00";  --  
tmp(170) := "000" & x"1" & '0' & x"01";  --  LDA $FLAG_INIBE_CONT
tmp(171) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(172) := "000" & x"7" & '0' & x"AF";  --  JEQ .incrementa_unidade
tmp(173) := "000" & x"A" & '0' & x"00";  --  RET
tmp(174) := "000" & x"0" & '0' & x"00";  --  
tmp(175) := "000" & x"0" & '0' & x"00";  --  incrementa_unidade:
tmp(176) := "000" & x"1" & '0' & x"02";  --  LDA $UNIDADE
tmp(177) := "000" & x"8" & '0' & x"0E";  --  CEQ $NOVE
tmp(178) := "000" & x"7" & '0' & x"B7";  --  JEQ .incrementa_dezena
tmp(179) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(180) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(181) := "000" & x"A" & '0' & x"00";  --  RET
tmp(182) := "000" & x"0" & '0' & x"00";  --  
tmp(183) := "000" & x"0" & '0' & x"00";  --  incrementa_dezena:
tmp(184) := "000" & x"1" & '0' & x"03";  --  LDA $DEZENA
tmp(185) := "000" & x"8" & '0' & x"11";  --  CEQ $CINCO
tmp(186) := "000" & x"7" & '0' & x"C1";  --  JEQ .incrementa_centena
tmp(187) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(188) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(189) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(190) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(191) := "000" & x"A" & '0' & x"00";  --  RET
tmp(192) := "000" & x"0" & '0' & x"00";  --  
tmp(193) := "000" & x"0" & '0' & x"00";  --  incrementa_centena:
tmp(194) := "000" & x"1" & '0' & x"04";  --  LDA $CENTENA
tmp(195) := "000" & x"8" & '0' & x"0E";  --  CEQ $NOVE
tmp(196) := "000" & x"7" & '0' & x"CC";  --  JEQ .incrementa_milhar
tmp(197) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(198) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(199) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(200) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(201) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(202) := "000" & x"A" & '0' & x"00";  --  RET
tmp(203) := "000" & x"0" & '0' & x"00";  --  
tmp(204) := "000" & x"0" & '0' & x"00";  --  incrementa_milhar:
tmp(205) := "000" & x"1" & '0' & x"05";  --  LDA $MILHAR
tmp(206) := "000" & x"8" & '0' & x"11";  --  CEQ $CINCO
tmp(207) := "000" & x"7" & '0' & x"D8";  --  JEQ .incrementa_dezena_milhar
tmp(208) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(209) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
tmp(210) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(211) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(212) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(213) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(214) := "000" & x"A" & '0' & x"00";  --  RET
tmp(215) := "000" & x"0" & '0' & x"00";  --  
tmp(216) := "000" & x"0" & '0' & x"00";  --  incrementa_dezena_milhar:
tmp(217) := "000" & x"1" & '0' & x"06";  --  LDA $DEZENA_MILHAR
tmp(218) := "000" & x"8" & '0' & x"12";  --  CEQ $TRES
tmp(219) := "000" & x"7" & '0' & x"E5";  --  JEQ .incrementa_centena_milhar
tmp(220) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(221) := "000" & x"5" & '0' & x"06";  --  STA $DEZENA_MILHAR
tmp(222) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(223) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(224) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(225) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(226) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
tmp(227) := "000" & x"A" & '0' & x"00";  --  RET
tmp(228) := "000" & x"0" & '0' & x"00";  --  
tmp(229) := "000" & x"0" & '0' & x"00";  --  incrementa_centena_milhar:
tmp(230) := "000" & x"1" & '0' & x"07";  --  LDA $CENTENA_MILHAR
tmp(231) := "000" & x"8" & '0' & x"10";  --  CEQ $DOIS
tmp(232) := "000" & x"7" & '0' & x"F3";  --  JEQ .zerar
tmp(233) := "000" & x"2" & '0' & x"0F";  --  SOMA $UM
tmp(234) := "000" & x"5" & '0' & x"07";  --  STA $CENTENA_MILHAR
tmp(235) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(236) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(237) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(238) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(239) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
tmp(240) := "000" & x"5" & '0' & x"06";  --  STA $DEZENA_MILHAR
tmp(241) := "000" & x"A" & '0' & x"00";  --  RET
tmp(242) := "000" & x"0" & '0' & x"00";  --  
tmp(243) := "000" & x"0" & '0' & x"00";  --  zerar:
tmp(244) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(245) := "000" & x"5" & '0' & x"02";  --  STA $UNIDADE
tmp(246) := "000" & x"5" & '0' & x"03";  --  STA $DEZENA
tmp(247) := "000" & x"5" & '0' & x"04";  --  STA $CENTENA
tmp(248) := "000" & x"5" & '0' & x"05";  --  STA $MILHAR
tmp(249) := "000" & x"5" & '0' & x"06";  --  STA $DEZENA_MILHAR
tmp(250) := "000" & x"5" & '0' & x"07";  --  STA $CENTENA_MILHAR
tmp(251) := "000" & x"A" & '0' & x"00";  --  RET
tmp(252) := "000" & x"0" & '0' & x"00";  --  
tmp(253) := "000" & x"0" & '0' & x"00";  --  limite:
tmp(254) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(255) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(256) := "000" & x"0" & '0' & x"00";  --  
tmp(257) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(258) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
tmp(259) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
tmp(260) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(261) := "000" & x"5" & '1' & x"23";  --  STA $HEX3
tmp(262) := "000" & x"5" & '1' & x"24";  --  STA $HEX4
tmp(263) := "000" & x"5" & '1' & x"25";  --  STA $HEX5
tmp(264) := "000" & x"0" & '0' & x"00";  --  
tmp(265) := "000" & x"0" & '0' & x"00";  --  ler_key1_und:
tmp(266) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(267) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(268) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(269) := "000" & x"7" & '1' & x"09";  --  JEQ .ler_key1_und
tmp(270) := "000" & x"0" & '0' & x"00";  --  
tmp(271) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(272) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(273) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(274) := "000" & x"5" & '0' & x"08";  --  STA $LIM_UNIDADE
tmp(275) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
tmp(276) := "000" & x"0" & '0' & x"00";  --  
tmp(277) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(278) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(279) := "000" & x"0" & '0' & x"00";  --  
tmp(280) := "000" & x"0" & '0' & x"00";  --  ler_key1_dez:
tmp(281) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(282) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(283) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(284) := "000" & x"7" & '1' & x"18";  --  JEQ .ler_key1_dez
tmp(285) := "000" & x"0" & '0' & x"00";  --  
tmp(286) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(287) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(288) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(289) := "000" & x"5" & '0' & x"09";  --  STA $LIM_DEZENA
tmp(290) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
tmp(291) := "000" & x"0" & '0' & x"00";  --  
tmp(292) := "000" & x"4" & '0' & x"03";  --  LDI $3
tmp(293) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(294) := "000" & x"0" & '0' & x"00";  --  
tmp(295) := "000" & x"0" & '0' & x"00";  --  ler_key1_cent:
tmp(296) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(297) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(298) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(299) := "000" & x"7" & '1' & x"27";  --  JEQ .ler_key1_cent
tmp(300) := "000" & x"0" & '0' & x"00";  --  
tmp(301) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(302) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(303) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(304) := "000" & x"5" & '0' & x"0A";  --  STA $LIM_CENTENA
tmp(305) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(306) := "000" & x"0" & '0' & x"00";  --  
tmp(307) := "000" & x"4" & '0' & x"07";  --  LDI $7
tmp(308) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(309) := "000" & x"0" & '0' & x"00";  --  
tmp(310) := "000" & x"0" & '0' & x"00";  --  ler_key1_mil:
tmp(311) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(312) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(313) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(314) := "000" & x"7" & '1' & x"36";  --  JEQ .ler_key1_mil
tmp(315) := "000" & x"0" & '0' & x"00";  --  
tmp(316) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(317) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(318) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(319) := "000" & x"5" & '0' & x"0B";  --  STA $LIM_MILHAR
tmp(320) := "000" & x"5" & '1' & x"23";  --  STA $HEX3
tmp(321) := "000" & x"0" & '0' & x"00";  --  
tmp(322) := "000" & x"4" & '0' & x"0F";  --  LDI $15
tmp(323) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(324) := "000" & x"0" & '0' & x"00";  --  
tmp(325) := "000" & x"0" & '0' & x"00";  --  ler_key1_dezmil:
tmp(326) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(327) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(328) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(329) := "000" & x"7" & '1' & x"45";  --  JEQ .ler_key1_dezmil
tmp(330) := "000" & x"0" & '0' & x"00";  --  
tmp(331) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(332) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(333) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(334) := "000" & x"5" & '0' & x"0C";  --  STA $LIM_DEZENA_MILHAR
tmp(335) := "000" & x"5" & '1' & x"24";  --  STA $HEX4
tmp(336) := "000" & x"0" & '0' & x"00";  --  
tmp(337) := "000" & x"4" & '0' & x"1F";  --  LDI $31
tmp(338) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(339) := "000" & x"0" & '0' & x"00";  --  
tmp(340) := "000" & x"0" & '0' & x"00";  --  ler_key1_centmil:
tmp(341) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(342) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(343) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(344) := "000" & x"7" & '1' & x"54";  --  JEQ .ler_key1_centmil
tmp(345) := "000" & x"0" & '0' & x"00";  --  
tmp(346) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(347) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(348) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(349) := "000" & x"5" & '0' & x"0D";  --  STA $LIM_CENTENA_MILHAR
tmp(350) := "000" & x"5" & '1' & x"25";  --  STA $HEX5
tmp(351) := "000" & x"0" & '0' & x"00";  --  
tmp(352) := "000" & x"4" & '0' & x"3F";  --  LDI $63
tmp(353) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(354) := "000" & x"0" & '0' & x"00";  --  
tmp(355) := "000" & x"0" & '0' & x"00";  --  ler_key1_after:
tmp(356) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(357) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(358) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(359) := "000" & x"7" & '1' & x"63";  --  JEQ .ler_key1_after
tmp(360) := "000" & x"0" & '0' & x"00";  --  
tmp(361) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(362) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(363) := "000" & x"0" & '0' & x"00";  --  
tmp(364) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(365) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(366) := "000" & x"0" & '0' & x"00";  --  
tmp(367) := "000" & x"1" & '0' & x"02";  --  LDA $UNIDADE
tmp(368) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
tmp(369) := "000" & x"0" & '0' & x"00";  --  
tmp(370) := "000" & x"1" & '0' & x"03";  --  LDA $DEZENA
tmp(371) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
tmp(372) := "000" & x"0" & '0' & x"00";  --  
tmp(373) := "000" & x"1" & '0' & x"04";  --  LDA $CENTENA
tmp(374) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(375) := "000" & x"0" & '0' & x"00";  --  
tmp(376) := "000" & x"1" & '0' & x"05";  --  LDA $MILHAR
tmp(377) := "000" & x"5" & '1' & x"23";  --  STA $HEX3
tmp(378) := "000" & x"0" & '0' & x"00";  --  
tmp(379) := "000" & x"1" & '0' & x"06";  --  LDA $DEZENA_MILHAR
tmp(380) := "000" & x"5" & '1' & x"24";  --  STA $HEX4
tmp(381) := "000" & x"0" & '0' & x"00";  --  
tmp(382) := "000" & x"1" & '0' & x"07";  --  LDA $CENTENA_MILHAR
tmp(383) := "000" & x"5" & '1' & x"25";  --  STA $HEX5
tmp(384) := "000" & x"0" & '0' & x"00";  --  
tmp(385) := "000" & x"A" & '0' & x"00";  --  RET

		
		
		return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;