library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDi : std_logic_vector(3 downto 0) := "1011";
  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  
   tmp(0) := "000" & x"4" & '0' & x"00";  --  LDI $0
  tmp(1) := "000" & x"5" & '0' & x"00";  --  STA $ZERO
  tmp(2) := "000" & x"0" & '0' & x"00";  --  
  tmp(3) := "000" & x"4" & '1' & x"FF";  --  LDI $511
  tmp(4) := "000" & x"0" & '0' & x"00";  --  
  tmp(5) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
  tmp(6) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
  tmp(7) := "000" & x"0" & '0' & x"00";  --  
  tmp(8) := "000" & x"4" & '0' & x"00";  --  LDI $0
  tmp(9) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
 tmp(10) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
 tmp(11) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
 tmp(12) := "000" & x"5" & '0' & x"01";  --  STA $LEDes
 tmp(13) := "000" & x"0" & '0' & x"00";  --  
 tmp(14) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
 tmp(15) := "000" & x"0" & '0' & x"00";  --  
 tmp(16) := "000" & x"5" & '0' & x"03";  --  STA $FLAG_INIBE_CONT
 tmp(17) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
 tmp(18) := "000" & x"5" & '1' & x"01";  --  STA $LEDR8
 tmp(19) := "000" & x"0" & '0' & x"00";  --  
 tmp(20) := "000" & x"5" & '0' & x"04";  --  STA $SEG
 tmp(21) := "000" & x"5" & '0' & x"05";  --  STA $MIN
 tmp(22) := "000" & x"5" & '0' & x"06";  --  STA $HR
 tmp(23) := "000" & x"5" & '0' & x"07";  --  STA $PM
 tmp(24) := "000" & x"0" & '0' & x"00";  --  
 tmp(25) := "000" & x"4" & '0' & x"01";  --  LDI $1
 tmp(26) := "000" & x"5" & '0' & x"08";  --  STA $UM
 tmp(27) := "000" & x"0" & '0' & x"00";  --  
 tmp(28) := "000" & x"0" & '0' & x"00";  --  
 tmp(29) := "000" & x"4" & '0' & x"3B";  --  LDI $59
 tmp(30) := "000" & x"5" & '0' & x"09";  --  STA $LIM_SEG
 tmp(31) := "000" & x"5" & '0' & x"0A";  --  STA $LIM_MIN
 tmp(32) := "000" & x"0" & '0' & x"00";  --  
 tmp(33) := "000" & x"0" & '0' & x"00";  --  
 tmp(34) := "000" & x"4" & '0' & x"17";  --  LDI $23
 tmp(35) := "000" & x"5" & '0' & x"0B";  --  STA $LIM_HR
 tmp(36) := "000" & x"0" & '0' & x"00";  --  
 tmp(37) := "000" & x"4" & '0' & x"0B";  --  LDI $11
 tmp(38) := "000" & x"5" & '0' & x"0C";  --  STA $LIM_HR_PM
 tmp(39) := "000" & x"0" & '0' & x"00";  --  
 tmp(40) := "000" & x"0" & '0' & x"00";  --  
 tmp(41) := "000" & x"0" & '0' & x"00";  --  main_loop:
 tmp(42) := "000" & x"0" & '0' & x"00";  --  
 tmp(43) := "000" & x"1" & '1' & x"60";  --  LDA $KEY0
 tmp(44) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(45) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(46) := "000" & x"7" & '0' & x"30";  --  JEQ .nao_leu_key0
 tmp(47) := "000" & x"9" & '0' & x"B3";  --  JSR .incrementa
 tmp(48) := "000" & x"0" & '0' & x"00";  --  nao_leu_key0:
 tmp(49) := "000" & x"0" & '0' & x"00";  --  
 tmp(50) := "000" & x"9" & '0' & x"41";  --  JSR .verifica_limite
 tmp(51) := "000" & x"0" & '0' & x"00";  --  
 tmp(52) := "000" & x"9" & '1' & x"09";  --  JSR .verifica_tipo
 tmp(53) := "000" & x"0" & '0' & x"00";  --  
 tmp(54) := "000" & x"1" & '0' & x"04";  --  LDA $SEG
 tmp(55) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
 tmp(56) := "000" & x"0" & '0' & x"00";  --  
 tmp(57) := "000" & x"1" & '0' & x"05";  --  LDA $MIN
 tmp(58) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
 tmp(59) := "000" & x"0" & '0' & x"00";  --  
 tmp(60) := "000" & x"0" & '0' & x"00";  --  
 tmp(61) := "000" & x"0" & '0' & x"00";  --  
 tmp(62) := "000" & x"0" & '0' & x"00";  --  
 tmp(63) := "000" & x"6" & '0' & x"29";  --  JMP .main_loop
 tmp(64) := "000" & x"0" & '0' & x"00";  --  
 tmp(65) := "000" & x"0" & '0' & x"00";  --  verifica_limite:
 tmp(66) := "000" & x"0" & '0' & x"00";  --  verifica_SEG:
 tmp(67) := "000" & x"1" & '0' & x"04";  --  LDA $SEG
 tmp(68) := "000" & x"8" & '0' & x"09";  --  CEQ $LIM_SEG
 tmp(69) := "000" & x"7" & '0' & x"48";  --  JEQ .verifica_MIN
 tmp(70) := "000" & x"A" & '0' & x"00";  --  RET
 tmp(71) := "000" & x"0" & '0' & x"00";  --  
 tmp(72) := "000" & x"0" & '0' & x"00";  --  verifica_MIN:
 tmp(73) := "000" & x"1" & '0' & x"05";  --  LDA $MIN
 tmp(74) := "000" & x"8" & '0' & x"0A";  --  CEQ $LIM_MIN
 tmp(75) := "000" & x"7" & '0' & x"4E";  --  JEQ .verifica_HR
 tmp(76) := "000" & x"A" & '0' & x"00";  --  RET
 tmp(77) := "000" & x"0" & '0' & x"00";  --  
 tmp(78) := "000" & x"0" & '0' & x"00";  --  verifica_HR:
 tmp(79) := "000" & x"1" & '0' & x"06";  --  LDA $HR
 tmp(80) := "000" & x"8" & '0' & x"0B";  --  CEQ $LIM_HR
 tmp(81) := "000" & x"7" & '0' & x"55";  --  JEQ .habilita_flag
 tmp(82) := "000" & x"A" & '0' & x"00";  --  RET
 tmp(83) := "000" & x"0" & '0' & x"00";  --  
 tmp(84) := "000" & x"0" & '0' & x"00";  --  
 tmp(85) := "000" & x"0" & '0' & x"00";  --  habilita_flag:
 tmp(86) := "000" & x"9" & '0' & x"5B";  --  JSR .dia_da_semana
 tmp(87) := "000" & x"0" & '0' & x"00";  --  
 tmp(88) := "000" & x"A" & '0' & x"00";  --  RET
 tmp(89) := "000" & x"0" & '0' & x"00";  --  
 tmp(90) := "000" & x"0" & '0' & x"00";  --  
 tmp(91) := "000" & x"0" & '0' & x"00";  --  dia_da_semana:
 tmp(92) := "000" & x"9" & '0' & x"5F";  --  JSR .calcula_dia
 tmp(93) := "000" & x"A" & '0' & x"00";  --  RET
 tmp(94) := "000" & x"0" & '0' & x"00";  --  
 tmp(95) := "000" & x"0" & '0' & x"00";  --  calcula_dia:
 tmp(96) := "000" & x"1" & '0' & x"0D";  --  LDA $DIA %8
 tmp(97) := "000" & x"2" & '0' & x"0E";  --  SOMA $UM %8
 tmp(98) := "000" & x"5" & '0' & x"0D";  --  STA $DIA %8
 tmp(99) := "000" & x"9" & '0' & x"6C";  --  JSR .verifica_dia
tmp(100) := "000" & x"A" & '0' & x"00";  --  RET
tmp(101) := "000" & x"0" & '0' & x"00";  --  
tmp(102) := "000" & x"0" & '0' & x"00";  --  rstdia:
tmp(103) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(104) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(105) := "000" & x"A" & '0' & x"00";  --  RET
tmp(106) := "000" & x"0" & '0' & x"00";  --  
tmp(107) := "000" & x"0" & '0' & x"00";  --  
tmp(108) := "000" & x"0" & '0' & x"00";  --  verifica_dia:
tmp(109) := "000" & x"1" & '0' & x"02";  --  LDA $DIA_N
tmp(110) := "000" & x"8" & '0' & x"02";  --  CEQ $2
tmp(111) := "000" & x"7" & '0' & x"7F";  --  JEQ .segunda
tmp(112) := "000" & x"8" & '0' & x"04";  --  CEQ $4
tmp(113) := "000" & x"7" & '0' & x"85";  --  JEQ .terca
tmp(114) := "000" & x"8" & '0' & x"08";  --  CEQ $8
tmp(115) := "000" & x"7" & '0' & x"8B";  --  JEQ .quarta
tmp(116) := "000" & x"8" & '0' & x"10";  --  CEQ $16
tmp(117) := "000" & x"7" & '0' & x"91";  --  JEQ .quinta
tmp(118) := "000" & x"8" & '0' & x"20";  --  CEQ $32
tmp(119) := "000" & x"7" & '0' & x"97";  --  JEQ .sexta
tmp(120) := "000" & x"8" & '0' & x"40";  --  CEQ $64
tmp(121) := "000" & x"7" & '0' & x"9D";  --  JEQ .sabado
tmp(122) := "000" & x"8" & '0' & x"80";  --  CEQ $128
tmp(123) := "000" & x"7" & '0' & x"A3";  --  JEQ .domingo
tmp(124) := "000" & x"9" & '0' & x"66";  --  JSR .rstdia
tmp(125) := "000" & x"A" & '0' & x"00";  --  RET
tmp(126) := "000" & x"0" & '0' & x"00";  --  
tmp(127) := "000" & x"0" & '0' & x"00";  --  segunda:
tmp(128) := "000" & x"4" & '0' & x"02";  --  LDI $2
tmp(129) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(130) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(131) := "000" & x"A" & '0' & x"00";  --  RET
tmp(132) := "000" & x"0" & '0' & x"00";  --  
tmp(133) := "000" & x"0" & '0' & x"00";  --  terca:
tmp(134) := "000" & x"4" & '0' & x"04";  --  LDI $4
tmp(135) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(136) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(137) := "000" & x"A" & '0' & x"00";  --  RET
tmp(138) := "000" & x"0" & '0' & x"00";  --  
tmp(139) := "000" & x"0" & '0' & x"00";  --  quarta:
tmp(140) := "000" & x"4" & '0' & x"08";  --  LDI $8
tmp(141) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(142) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(143) := "000" & x"A" & '0' & x"00";  --  RET
tmp(144) := "000" & x"0" & '0' & x"00";  --  
tmp(145) := "000" & x"0" & '0' & x"00";  --  quinta:
tmp(146) := "000" & x"4" & '0' & x"10";  --  LDI $16
tmp(147) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(148) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(149) := "000" & x"A" & '0' & x"00";  --  RET
tmp(150) := "000" & x"0" & '0' & x"00";  --  
tmp(151) := "000" & x"0" & '0' & x"00";  --  sexta:
tmp(152) := "000" & x"4" & '0' & x"20";  --  LDI $32
tmp(153) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(154) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(155) := "000" & x"A" & '0' & x"00";  --  RET
tmp(156) := "000" & x"0" & '0' & x"00";  --  
tmp(157) := "000" & x"0" & '0' & x"00";  --  sabado:
tmp(158) := "000" & x"4" & '0' & x"40";  --  LDI $64
tmp(159) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(160) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(161) := "000" & x"A" & '0' & x"00";  --  RET
tmp(162) := "000" & x"0" & '0' & x"00";  --  
tmp(163) := "000" & x"0" & '0' & x"00";  --  domingo:
tmp(164) := "000" & x"4" & '0' & x"80";  --  LDI $128
tmp(165) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(166) := "000" & x"5" & '0' & x"02";  --  STA $DIA_N
tmp(167) := "000" & x"A" & '0' & x"00";  --  RET
tmp(168) := "000" & x"0" & '0' & x"00";  --  
tmp(169) := "000" & x"0" & '0' & x"00";  --  
tmp(170) := "000" & x"0" & '0' & x"00";  --  
tmp(171) := "000" & x"0" & '0' & x"00";  --  reset:
tmp(172) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(173) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(174) := "000" & x"5" & '0' & x"05";  --  STA $MIN
tmp(175) := "000" & x"5" & '0' & x"06";  --  STA $HR
tmp(176) := "000" & x"5" & '0' & x"07";  --  STA $PM
tmp(177) := "000" & x"A" & '0' & x"00";  --  RET
tmp(178) := "000" & x"0" & '0' & x"00";  --  
tmp(179) := "000" & x"0" & '0' & x"00";  --  incrementa:
tmp(180) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(181) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
tmp(182) := "000" & x"0" & '0' & x"00";  --  
tmp(183) := "000" & x"1" & '0' & x"03";  --  LDA $FLAG_INIBE_CONT
tmp(184) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(185) := "000" & x"7" & '0' & x"BC";  --  JEQ .incrementa_SEG
tmp(186) := "000" & x"A" & '0' & x"00";  --  RET
tmp(187) := "000" & x"0" & '0' & x"00";  --  
tmp(188) := "000" & x"0" & '0' & x"00";  --  incrementa_SEG:
tmp(189) := "000" & x"1" & '0' & x"04";  --  LDA $SEG
tmp(190) := "000" & x"8" & '0' & x"09";  --  CEQ $LIM_SEG
tmp(191) := "000" & x"7" & '0' & x"C4";  --  JEQ .incrementa_MIN
tmp(192) := "000" & x"2" & '0' & x"08";  --  SOMA $UM
tmp(193) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(194) := "000" & x"A" & '0' & x"00";  --  RET
tmp(195) := "000" & x"0" & '0' & x"00";  --  
tmp(196) := "000" & x"0" & '0' & x"00";  --  incrementa_MIN:
tmp(197) := "000" & x"1" & '0' & x"05";  --  LDA $MIN
tmp(198) := "000" & x"8" & '0' & x"0A";  --  CEQ $LIM_MIN
tmp(199) := "000" & x"7" & '0' & x"CE";  --  JEQ .incrementa_HR
tmp(200) := "000" & x"2" & '0' & x"08";  --  SOMA $UM
tmp(201) := "000" & x"5" & '0' & x"05";  --  STA $MIN
tmp(202) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(203) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(204) := "000" & x"A" & '0' & x"00";  --  RET
tmp(205) := "000" & x"0" & '0' & x"00";  --  
tmp(206) := "000" & x"0" & '0' & x"00";  --  incrementa_HR:
tmp(207) := "000" & x"1" & '0' & x"0F";  --  LDA $FLAG_PM
tmp(208) := "000" & x"8" & '0' & x"08";  --  CEQ $UM
tmp(209) := "000" & x"7" & '0' & x"DC";  --  JEQ .incrementa_HR_PM
tmp(210) := "000" & x"1" & '0' & x"06";  --  LDA $HR
tmp(211) := "000" & x"8" & '0' & x"0B";  --  CEQ $LIM_HR
tmp(212) := "000" & x"7" & '0' & x"E7";  --  JEQ .zerar
tmp(213) := "000" & x"2" & '0' & x"08";  --  SOMA $UM
tmp(214) := "000" & x"5" & '0' & x"06";  --  STA $HR
tmp(215) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(216) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(217) := "000" & x"5" & '0' & x"05";  --  STA $MIN
tmp(218) := "000" & x"A" & '0' & x"00";  --  RET
tmp(219) := "000" & x"0" & '0' & x"00";  --  
tmp(220) := "000" & x"0" & '0' & x"00";  --  incrementa_HR_PM:
tmp(221) := "000" & x"1" & '0' & x"07";  --  LDA $PM
tmp(222) := "000" & x"8" & '0' & x"0C";  --  CEQ $LIM_HR_PM
tmp(223) := "000" & x"7" & '0' & x"E7";  --  JEQ .zerar
tmp(224) := "000" & x"2" & '0' & x"08";  --  SOMA $UM
tmp(225) := "000" & x"5" & '0' & x"07";  --  STA $PM
tmp(226) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(227) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(228) := "000" & x"5" & '0' & x"05";  --  STA $MIN
tmp(229) := "000" & x"A" & '0' & x"00";  --  RET
tmp(230) := "000" & x"0" & '0' & x"00";  --  
tmp(231) := "000" & x"0" & '0' & x"00";  --  zerar:
tmp(232) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(233) := "000" & x"5" & '0' & x"04";  --  STA $SEG
tmp(234) := "000" & x"5" & '0' & x"05";  --  STA $MIN
tmp(235) := "000" & x"5" & '0' & x"06";  --  STA $HR
tmp(236) := "000" & x"5" & '0' & x"07";  --  STA $PM
tmp(237) := "000" & x"1" & '0' & x"0F";  --  LDA $FLAG_PM
tmp(238) := "000" & x"8" & '0' & x"08";  --  CEQ $UM
tmp(239) := "000" & x"7" & '0' & x"F6";  --  JEQ .ativa_led_PM
tmp(240) := "000" & x"1" & '0' & x"01";  --  LDA $LEDes
tmp(241) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(242) := "000" & x"5" & '0' & x"01";  --  STA $LEDes
tmp(243) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(244) := "000" & x"A" & '0' & x"00";  --  RET
tmp(245) := "000" & x"0" & '0' & x"00";  --  
tmp(246) := "000" & x"0" & '0' & x"00";  --  ativa_led_PM:
tmp(247) := "000" & x"9" & '0' & x"FA";  --  JSR .logica_PM
tmp(248) := "000" & x"A" & '0' & x"00";  --  RET
tmp(249) := "000" & x"0" & '0' & x"00";  --  
tmp(250) := "000" & x"0" & '0' & x"00";  --  logica_PM:
tmp(251) := "000" & x"1" & '0' & x"01";  --  LDA $LEDes
tmp(252) := "000" & x"8" & '0' & x"01";  --  CEQ $1
tmp(253) := "000" & x"7" & '1' & x"03";  --  JEQ .desativa_PM
tmp(254) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(255) := "000" & x"5" & '0' & x"01";  --  STA $LEDes
tmp(256) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(257) := "000" & x"A" & '0' & x"00";  --  RET
tmp(258) := "000" & x"0" & '0' & x"00";  --  
tmp(259) := "000" & x"0" & '0' & x"00";  --  desativa_PM:
tmp(260) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(261) := "000" & x"5" & '0' & x"01";  --  STA $LEDes
tmp(262) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(263) := "000" & x"A" & '0' & x"00";  --  RET
tmp(264) := "000" & x"0" & '0' & x"00";  --  
tmp(265) := "000" & x"0" & '0' & x"00";  --  verifica_tipo:
tmp(266) := "000" & x"1" & '1' & x"41";  --  LDA $SW8
tmp(267) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(268) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(269) := "000" & x"0" & '0' & x"00";  --  
tmp(270) := "000" & x"7" & '1' & x"16";  --  JEQ .ativa_PM
tmp(271) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(272) := "000" & x"5" & '0' & x"0F";  --  STA $FLAG_PM
tmp(273) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(274) := "000" & x"1" & '0' & x"06";  --  LDA $HR
tmp(275) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(276) := "000" & x"A" & '0' & x"00";  --  RET
tmp(277) := "000" & x"0" & '0' & x"00";  --  
tmp(278) := "000" & x"0" & '0' & x"00";  --  ativa_PM:
tmp(279) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(280) := "000" & x"5" & '0' & x"0F";  --  STA $FLAG_PM
tmp(281) := "000" & x"1" & '0' & x"07";  --  LDA $PM
tmp(282) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(283) := "000" & x"A" & '0' & x"00";  --  RET



		
		return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;