library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDi : std_logic_vector(3 downto 0) := "1011";
  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  
  tmp(0) := "000" & x"4" & '0' & x"00";  --  LDI $0
  tmp(1) := "000" & x"5" & '0' & x"00";  --  STA $ZERO
  tmp(2) := "000" & x"0" & '0' & x"00";  --  
  tmp(3) := "000" & x"4" & '0' & x"01";  --  LDI $1
  tmp(4) := "000" & x"5" & '0' & x"01";  --  STA $UM
  tmp(5) := "000" & x"0" & '0' & x"00";  --  
  tmp(6) := "001" & x"4" & '1' & x"FF";  --  LDI $511 %1
  tmp(7) := "000" & x"5" & '0' & x"02";  --  STA $CLR_KEY0 %1
  tmp(8) := "000" & x"5" & '0' & x"03";  --  STA $CLR_KEY1 %1
  tmp(9) := "000" & x"5" & '0' & x"04";  --  STA $CLR_KEY2 %1
 tmp(10) := "000" & x"5" & '0' & x"05";  --  STA $CLR_KEY3 %1
 tmp(11) := "000" & x"0" & '0' & x"00";  --  
 tmp(12) := "000" & x"4" & '0' & x"00";  --  LDI $0
 tmp(13) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
 tmp(14) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
 tmp(15) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
 tmp(16) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
 tmp(17) := "000" & x"0" & '0' & x"00";  --  
 tmp(18) := "000" & x"5" & '0' & x"06";  --  STA $FLAG_DESPERTADOR
 tmp(19) := "000" & x"5" & '1' & x"02";  --  STA $LEDR9
 tmp(20) := "000" & x"5" & '1' & x"01";  --  STA $LEDR8
 tmp(21) := "000" & x"0" & '0' & x"00";  --  
 tmp(22) := "000" & x"5" & '0' & x"07";  --  STA $SEG
 tmp(23) := "000" & x"5" & '0' & x"08";  --  STA $MIN
 tmp(24) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
 tmp(25) := "000" & x"5" & '0' & x"0A";  --  STA $HR_12
 tmp(26) := "000" & x"0" & '0' & x"00";  --  
 tmp(27) := "000" & x"4" & '0' & x"3B";  --  LDI $59
 tmp(28) := "000" & x"5" & '0' & x"0B";  --  STA $LIM_SEG
 tmp(29) := "000" & x"5" & '0' & x"0C";  --  STA $LIM_MIN
 tmp(30) := "000" & x"0" & '0' & x"00";  --  
 tmp(31) := "000" & x"4" & '0' & x"17";  --  LDI $23
 tmp(32) := "000" & x"5" & '0' & x"0D";  --  STA $LIM_HR_24
 tmp(33) := "000" & x"0" & '0' & x"00";  --  
 tmp(34) := "000" & x"4" & '0' & x"0B";  --  LDI $11
 tmp(35) := "000" & x"5" & '0' & x"0E";  --  STA $LIM_HR_12
 tmp(36) := "000" & x"0" & '0' & x"00";  --  
 tmp(37) := "000" & x"4" & '0' & x"00";  --  LDI $0
 tmp(38) := "000" & x"5" & '0' & x"0F";  --  STA $DESP_HORAS
 tmp(39) := "000" & x"5" & '0' & x"10";  --  STA $DESP_MINUTOS
 tmp(40) := "000" & x"4" & '0' & x"2D";  --  LDI $45
 tmp(41) := "000" & x"5" & '0' & x"11";  --  STA $DESP_SEGUNDOS
 tmp(42) := "000" & x"0" & '0' & x"00";  --  
 tmp(43) := "000" & x"0" & '0' & x"00";  --  volta_main_loop:
 tmp(44) := "000" & x"4" & '1' & x"FF";  --  LDI $511
 tmp(45) := "000" & x"5" & '1' & x"FD";  --  STA $CLR_KEY2
 tmp(46) := "000" & x"0" & '0' & x"00";  --  
 tmp(47) := "000" & x"0" & '0' & x"00";  --  main_loop:
 tmp(48) := "000" & x"1" & '1' & x"60";  --  LDA $KEY0
 tmp(49) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(50) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(51) := "000" & x"7" & '0' & x"41";  --  JEQ .nao_leu_key0
 tmp(52) := "000" & x"1" & '1' & x"41";  --  LDA $SW8
 tmp(53) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(54) := "000" & x"8" & '0' & x"01";  --  CEQ $1
 tmp(55) := "000" & x"7" & '0' & x"39";  --  JEQ .not_inverted
 tmp(56) := "000" & x"9" & '1' & x"28";  --  JSR .incrementa_segundos
 tmp(57) := "000" & x"0" & '0' & x"00";  --  not_inverted:
 tmp(58) := "000" & x"0" & '0' & x"00";  --  
 tmp(59) := "000" & x"1" & '1' & x"41";  --  LDA $SW8
 tmp(60) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(61) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(62) := "000" & x"7" & '0' & x"40";  --  JEQ .inverted
 tmp(63) := "000" & x"9" & '0' & x"FF";  --  JSR .decrementa_segundos
 tmp(64) := "000" & x"0" & '0' & x"00";  --  inverted:
 tmp(65) := "000" & x"0" & '0' & x"00";  --  nao_leu_key0:
 tmp(66) := "000" & x"0" & '0' & x"00";  --  
 tmp(67) := "000" & x"1" & '1' & x"62";  --  LDA $KEY2
 tmp(68) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(69) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(70) := "000" & x"7" & '0' & x"48";  --  JEQ .nao_leu_key2
 tmp(71) := "000" & x"9" & '0' & x"58";  --  JSR .define_segundos_horario
 tmp(72) := "000" & x"0" & '0' & x"00";  --  nao_leu_key2:
 tmp(73) := "000" & x"0" & '0' & x"00";  --  
 tmp(74) := "000" & x"1" & '1' & x"64";  --  LDA $FPGA_RESET
 tmp(75) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(76) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(77) := "000" & x"7" & '0' & x"50";  --  JEQ .nao_leu_reset
 tmp(78) := "000" & x"4" & '0' & x"00";  --  LDI $0
 tmp(79) := "000" & x"5" & '0' & x"06";  --  STA $FLAG_DESPERTADOR
 tmp(80) := "000" & x"0" & '0' & x"00";  --  nao_leu_reset:
 tmp(81) := "000" & x"0" & '0' & x"00";  --  
 tmp(82) := "000" & x"9" & '1' & x"51";  --  JSR .atualiza_display_horario
 tmp(83) := "000" & x"0" & '0' & x"00";  --  
 tmp(84) := "000" & x"9" & '0' & x"D6";  --  JSR .verifica_flag_despertador
 tmp(85) := "000" & x"0" & '0' & x"00";  --  
 tmp(86) := "000" & x"6" & '0' & x"2F";  --  JMP .main_loop
 tmp(87) := "000" & x"0" & '0' & x"00";  --  
 tmp(88) := "000" & x"0" & '0' & x"00";  --  define_segundos_horario:
 tmp(89) := "000" & x"4" & '1' & x"FF";  --  LDI $511
 tmp(90) := "000" & x"5" & '1' & x"FD";  --  STA $CLR_KEY2
 tmp(91) := "000" & x"0" & '0' & x"00";  --  
 tmp(92) := "000" & x"0" & '0' & x"00";  --  loop_define_segundos_horario:
 tmp(93) := "000" & x"4" & '0' & x"03";  --  LDI $3
 tmp(94) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
 tmp(95) := "000" & x"0" & '0' & x"00";  --  
 tmp(96) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
 tmp(97) := "000" & x"B" & '0' & x"01";  --  ANDI $1
 tmp(98) := "000" & x"8" & '0' & x"00";  --  CEQ $0
 tmp(99) := "000" & x"7" & '0' & x"65";  --  JEQ .nao_leu_key1_def_hor
tmp(100) := "000" & x"9" & '0' & x"A6";  --  JSR .def_horario_incrementa_segundos
tmp(101) := "000" & x"0" & '0' & x"00";  --  nao_leu_key1_def_hor:
tmp(102) := "000" & x"0" & '0' & x"00";  --  
tmp(103) := "000" & x"1" & '1' & x"62";  --  LDA $KEY2
tmp(104) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(105) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(106) := "000" & x"7" & '0' & x"6C";  --  JEQ .nao_leu_key2_def_hor
tmp(107) := "000" & x"9" & '0' & x"72";  --  JSR .define_minutos_horario
tmp(108) := "000" & x"0" & '0' & x"00";  --  nao_leu_key2_def_hor:
tmp(109) := "000" & x"0" & '0' & x"00";  --  
tmp(110) := "000" & x"9" & '1' & x"51";  --  JSR .atualiza_display_horario
tmp(111) := "000" & x"0" & '0' & x"00";  --  
tmp(112) := "000" & x"6" & '0' & x"5C";  --  JMP .loop_define_segundos_horario
tmp(113) := "000" & x"0" & '0' & x"00";  --  
tmp(114) := "000" & x"0" & '0' & x"00";  --  define_minutos_horario:
tmp(115) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(116) := "000" & x"5" & '1' & x"FD";  --  STA $CLR_KEY2
tmp(117) := "000" & x"0" & '0' & x"00";  --  
tmp(118) := "000" & x"0" & '0' & x"00";  --  loop_define_minutos_horario:
tmp(119) := "000" & x"4" & '0' & x"18";  --  LDI $24
tmp(120) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(121) := "000" & x"0" & '0' & x"00";  --  
tmp(122) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(123) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(124) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(125) := "000" & x"7" & '0' & x"7F";  --  JEQ .nao_leu_key1_def_min
tmp(126) := "000" & x"9" & '0' & x"B6";  --  JSR .def_horario_incrementa_minutos
tmp(127) := "000" & x"0" & '0' & x"00";  --  nao_leu_key1_def_min:
tmp(128) := "000" & x"0" & '0' & x"00";  --  
tmp(129) := "000" & x"1" & '1' & x"62";  --  LDA $KEY2
tmp(130) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(131) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(132) := "000" & x"7" & '0' & x"86";  --  JEQ .nao_leu_key2_def_min
tmp(133) := "000" & x"9" & '0' & x"8C";  --  JSR .define_horas_horario
tmp(134) := "000" & x"0" & '0' & x"00";  --  nao_leu_key2_def_min:
tmp(135) := "000" & x"0" & '0' & x"00";  --  
tmp(136) := "000" & x"9" & '1' & x"51";  --  JSR .atualiza_display_horario
tmp(137) := "000" & x"0" & '0' & x"00";  --  
tmp(138) := "000" & x"6" & '0' & x"76";  --  JMP .loop_define_minutos_horario
tmp(139) := "000" & x"0" & '0' & x"00";  --  
tmp(140) := "000" & x"0" & '0' & x"00";  --  define_horas_horario:
tmp(141) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(142) := "000" & x"5" & '1' & x"FD";  --  STA $CLR_KEY2
tmp(143) := "000" & x"0" & '0' & x"00";  --  
tmp(144) := "000" & x"0" & '0' & x"00";  --  loop_define_horas_horario:
tmp(145) := "000" & x"4" & '0' & x"C0";  --  LDI $192
tmp(146) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(147) := "000" & x"0" & '0' & x"00";  --  
tmp(148) := "000" & x"1" & '1' & x"61";  --  LDA $KEY1
tmp(149) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(150) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(151) := "000" & x"7" & '0' & x"99";  --  JEQ .nao_leu_key1_def_hr
tmp(152) := "000" & x"9" & '0' & x"C6";  --  JSR .def_horario_incrementa_horas
tmp(153) := "000" & x"0" & '0' & x"00";  --  nao_leu_key1_def_hr:
tmp(154) := "000" & x"0" & '0' & x"00";  --  
tmp(155) := "000" & x"1" & '1' & x"62";  --  LDA $KEY2
tmp(156) := "000" & x"B" & '0' & x"01";  --  ANDI $1
tmp(157) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(158) := "000" & x"7" & '0' & x"A0";  --  JEQ .nao_leu_key2_def_hr
tmp(159) := "000" & x"6" & '0' & x"2B";  --  JMP .volta_main_loop
tmp(160) := "000" & x"0" & '0' & x"00";  --  nao_leu_key2_def_hr:
tmp(161) := "000" & x"0" & '0' & x"00";  --  
tmp(162) := "000" & x"9" & '1' & x"51";  --  JSR .atualiza_display_horario
tmp(163) := "000" & x"0" & '0' & x"00";  --  
tmp(164) := "000" & x"6" & '0' & x"90";  --  JMP .loop_define_horas_horario
tmp(165) := "000" & x"0" & '0' & x"00";  --  
tmp(166) := "000" & x"0" & '0' & x"00";  --  def_horario_incrementa_segundos:
tmp(167) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(168) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(169) := "000" & x"0" & '0' & x"00";  --  
tmp(170) := "000" & x"1" & '0' & x"07";  --  LDA $SEG
tmp(171) := "000" & x"8" & '0' & x"0B";  --  CEQ $LIM_SEG
tmp(172) := "000" & x"7" & '0' & x"B1";  --  JEQ .def_horario_zera_segundos
tmp(173) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(174) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(175) := "000" & x"A" & '0' & x"00";  --  RET
tmp(176) := "000" & x"0" & '0' & x"00";  --  
tmp(177) := "000" & x"0" & '0' & x"00";  --  def_horario_zera_segundos:
tmp(178) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(179) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(180) := "000" & x"A" & '0' & x"00";  --  RET
tmp(181) := "000" & x"0" & '0' & x"00";  --  
tmp(182) := "000" & x"0" & '0' & x"00";  --  def_horario_incrementa_minutos:
tmp(183) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(184) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(185) := "000" & x"0" & '0' & x"00";  --  
tmp(186) := "000" & x"1" & '0' & x"08";  --  LDA $MIN
tmp(187) := "000" & x"8" & '0' & x"0C";  --  CEQ $LIM_MIN
tmp(188) := "000" & x"7" & '0' & x"C1";  --  JEQ .def_horario_zera_minutos
tmp(189) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(190) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(191) := "000" & x"A" & '0' & x"00";  --  RET
tmp(192) := "000" & x"0" & '0' & x"00";  --  
tmp(193) := "000" & x"0" & '0' & x"00";  --  def_horario_zera_minutos:
tmp(194) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(195) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(196) := "000" & x"A" & '0' & x"00";  --  RET
tmp(197) := "000" & x"0" & '0' & x"00";  --  
tmp(198) := "000" & x"0" & '0' & x"00";  --  def_horario_incrementa_horas:
tmp(199) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(200) := "000" & x"5" & '1' & x"FE";  --  STA $CLR_KEY1
tmp(201) := "000" & x"0" & '0' & x"00";  --  
tmp(202) := "000" & x"1" & '0' & x"09";  --  LDA $HR_24
tmp(203) := "000" & x"8" & '0' & x"0D";  --  CEQ $LIM_HR_24
tmp(204) := "000" & x"7" & '0' & x"D1";  --  JEQ .def_horario_zera_horas
tmp(205) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(206) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
tmp(207) := "000" & x"A" & '0' & x"00";  --  RET
tmp(208) := "000" & x"0" & '0' & x"00";  --  
tmp(209) := "000" & x"0" & '0' & x"00";  --  def_horario_zera_horas:
tmp(210) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(211) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
tmp(212) := "000" & x"A" & '0' & x"00";  --  RET
tmp(213) := "000" & x"0" & '0' & x"00";  --  
tmp(214) := "000" & x"0" & '0' & x"00";  --  verifica_flag_despertador:
tmp(215) := "000" & x"1" & '0' & x"06";  --  LDA $FLAG_DESPERTADOR
tmp(216) := "000" & x"8" & '0' & x"00";  --  CEQ $0
tmp(217) := "000" & x"7" & '0' & x"E2";  --  JEQ .apaga_leds
tmp(218) := "000" & x"9" & '0' & x"DD";  --  JSR .acende_leds
tmp(219) := "000" & x"A" & '0' & x"00";  --  RET
tmp(220) := "000" & x"0" & '0' & x"00";  --  
tmp(221) := "000" & x"0" & '0' & x"00";  --  acende_leds:
tmp(222) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(223) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(224) := "000" & x"A" & '0' & x"00";  --  RET
tmp(225) := "000" & x"0" & '0' & x"00";  --  
tmp(226) := "000" & x"0" & '0' & x"00";  --  apaga_leds:
tmp(227) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(228) := "000" & x"5" & '1' & x"00";  --  STA $LEDS
tmp(229) := "000" & x"A" & '0' & x"00";  --  RET
tmp(230) := "000" & x"0" & '0' & x"00";  --  
tmp(231) := "000" & x"0" & '0' & x"00";  --  verifica_despertador:
tmp(232) := "000" & x"1" & '0' & x"07";  --  LDA $SEG
tmp(233) := "000" & x"8" & '0' & x"11";  --  CEQ $DESP_SEGUNDOS
tmp(234) := "000" & x"7" & '0' & x"ED";  --  JEQ .verifica_minutos_despertador
tmp(235) := "000" & x"A" & '0' & x"00";  --  RET
tmp(236) := "000" & x"0" & '0' & x"00";  --  
tmp(237) := "000" & x"0" & '0' & x"00";  --  verifica_minutos_despertador:
tmp(238) := "000" & x"1" & '0' & x"08";  --  LDA $MIN
tmp(239) := "000" & x"8" & '0' & x"10";  --  CEQ $DESP_MINUTOS
tmp(240) := "000" & x"7" & '0' & x"F3";  --  JEQ .verifica_horas_despertador
tmp(241) := "000" & x"A" & '0' & x"00";  --  RET
tmp(242) := "000" & x"0" & '0' & x"00";  --  
tmp(243) := "000" & x"0" & '0' & x"00";  --  verifica_horas_despertador:
tmp(244) := "000" & x"1" & '1' & x"40";  --  LDA $SWS
tmp(245) := "000" & x"B" & '0' & x"7F";  --  ANDI $127
tmp(246) := "000" & x"8" & '0' & x"09";  --  CEQ $HR_24
tmp(247) := "000" & x"7" & '0' & x"FA";  --  JEQ .despertou
tmp(248) := "000" & x"A" & '0' & x"00";  --  RET
tmp(249) := "000" & x"0" & '0' & x"00";  --  
tmp(250) := "000" & x"0" & '0' & x"00";  --  despertou:
tmp(251) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(252) := "000" & x"5" & '0' & x"06";  --  STA $FLAG_DESPERTADOR
tmp(253) := "000" & x"A" & '0' & x"00";  --  RET
tmp(254) := "000" & x"0" & '0' & x"00";  --  
tmp(255) := "000" & x"0" & '0' & x"00";  --  decrementa_segundos:
tmp(256) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(257) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
tmp(258) := "000" & x"0" & '0' & x"00";  --  
tmp(259) := "000" & x"4" & '0' & x"00";  --  LDI $0
tmp(260) := "000" & x"5" & '0' & x"06";  --  STA $FLAG_DESPERTADOR
tmp(261) := "000" & x"0" & '0' & x"00";  --  
tmp(262) := "000" & x"1" & '0' & x"07";  --  LDA $SEG
tmp(263) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(264) := "000" & x"7" & '1' & x"0D";  --  JEQ .decrementa_minutos
tmp(265) := "000" & x"3" & '0' & x"01";  --  SUB $UM
tmp(266) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(267) := "000" & x"A" & '0' & x"00";  --  RET
tmp(268) := "000" & x"0" & '0' & x"00";  --  
tmp(269) := "000" & x"0" & '0' & x"00";  --  decrementa_minutos:
tmp(270) := "000" & x"1" & '0' & x"08";  --  LDA $MIN
tmp(271) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(272) := "000" & x"7" & '1' & x"17";  --  JEQ .decrementa_horas
tmp(273) := "000" & x"3" & '0' & x"01";  --  SUB $UM
tmp(274) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(275) := "000" & x"1" & '0' & x"0B";  --  LDA $LIM_SEG
tmp(276) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(277) := "000" & x"A" & '0' & x"00";  --  RET
tmp(278) := "000" & x"0" & '0' & x"00";  --  
tmp(279) := "000" & x"0" & '0' & x"00";  --  decrementa_horas:
tmp(280) := "000" & x"1" & '0' & x"09";  --  LDA $HR_24
tmp(281) := "000" & x"8" & '0' & x"00";  --  CEQ $ZERO
tmp(282) := "000" & x"7" & '1' & x"23";  --  JEQ .down_zera
tmp(283) := "000" & x"3" & '0' & x"01";  --  SUB $UM
tmp(284) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
tmp(285) := "000" & x"1" & '0' & x"0C";  --  LDA $LIM_MIN
tmp(286) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(287) := "000" & x"1" & '0' & x"0B";  --  LDA $LIM_SEG
tmp(288) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(289) := "000" & x"A" & '0' & x"00";  --  RET
tmp(290) := "000" & x"0" & '0' & x"00";  --  
tmp(291) := "000" & x"0" & '0' & x"00";  --  down_zera:
tmp(292) := "000" & x"4" & '0' & x"01";  --  LDI $1
tmp(293) := "000" & x"5" & '0' & x"06";  --  STA $FLAG_DESPERTADOR
tmp(294) := "000" & x"A" & '0' & x"00";  --  RET
tmp(295) := "000" & x"0" & '0' & x"00";  --  
tmp(296) := "000" & x"0" & '0' & x"00";  --  incrementa_segundos:
tmp(297) := "000" & x"4" & '1' & x"FF";  --  LDI $511
tmp(298) := "000" & x"5" & '1' & x"FF";  --  STA $CLR_KEY0
tmp(299) := "000" & x"0" & '0' & x"00";  --  
tmp(300) := "000" & x"9" & '0' & x"E7";  --  JSR .verifica_despertador
tmp(301) := "000" & x"0" & '0' & x"00";  --  
tmp(302) := "000" & x"1" & '0' & x"07";  --  LDA $SEG
tmp(303) := "000" & x"8" & '0' & x"0B";  --  CEQ $LIM_SEG
tmp(304) := "000" & x"7" & '1' & x"35";  --  JEQ .incrementa_minutos
tmp(305) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(306) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(307) := "000" & x"A" & '0' & x"00";  --  RET
tmp(308) := "000" & x"0" & '0' & x"00";  --  
tmp(309) := "000" & x"0" & '0' & x"00";  --  incrementa_minutos:
tmp(310) := "000" & x"1" & '0' & x"08";  --  LDA $MIN
tmp(311) := "000" & x"8" & '0' & x"0C";  --  CEQ $LIM_MIN
tmp(312) := "000" & x"7" & '1' & x"3F";  --  JEQ .incrementa_horas
tmp(313) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(314) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(315) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(316) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(317) := "000" & x"A" & '0' & x"00";  --  RET
tmp(318) := "000" & x"0" & '0' & x"00";  --  
tmp(319) := "000" & x"0" & '0' & x"00";  --  incrementa_horas:
tmp(320) := "000" & x"1" & '0' & x"09";  --  LDA $HR_24
tmp(321) := "000" & x"8" & '0' & x"0D";  --  CEQ $LIM_HR_24
tmp(322) := "000" & x"7" & '1' & x"4A";  --  JEQ .zera
tmp(323) := "000" & x"2" & '0' & x"01";  --  SOMA $UM
tmp(324) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
tmp(325) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(326) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(327) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(328) := "000" & x"A" & '0' & x"00";  --  RET
tmp(329) := "000" & x"0" & '0' & x"00";  --  
tmp(330) := "000" & x"0" & '0' & x"00";  --  zera:
tmp(331) := "000" & x"1" & '0' & x"00";  --  LDA $ZERO
tmp(332) := "000" & x"5" & '0' & x"09";  --  STA $HR_24
tmp(333) := "000" & x"5" & '0' & x"08";  --  STA $MIN
tmp(334) := "000" & x"5" & '0' & x"07";  --  STA $SEG
tmp(335) := "000" & x"A" & '0' & x"00";  --  RET
tmp(336) := "000" & x"0" & '0' & x"00";  --  
tmp(337) := "000" & x"0" & '0' & x"00";  --  atualiza_display_horario:
tmp(338) := "000" & x"1" & '0' & x"07";  --  LDA $SEG
tmp(339) := "000" & x"5" & '1' & x"20";  --  STA $HEX0
tmp(340) := "000" & x"0" & '0' & x"00";  --  
tmp(341) := "000" & x"1" & '0' & x"08";  --  LDA $MIN
tmp(342) := "000" & x"5" & '1' & x"21";  --  STA $HEX1
tmp(343) := "000" & x"0" & '0' & x"00";  --  
tmp(344) := "000" & x"1" & '0' & x"09";  --  LDA $HR_24
tmp(345) := "000" & x"5" & '1' & x"22";  --  STA $HEX2
tmp(346) := "000" & x"A" & '0' & x"00";  --  RET
		return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;